module external_mod(input[15:0] x, output[15:0] __output);
    assign __output = x+1;
endmodule
